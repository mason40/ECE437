`include "cpu_types_pkg.vh"

import cpu_types_pkg::*;

// module declaration
module alu (
